library IEEE;
use IEEE.std_logic_1164.all;

use work.my_components.all;

